`ifndef PARAMETER_H
DEFINE PARAMETER_H

`define b_width       16
`define i_width       8
`define mem_size      65536
`define ram_size      4095

`endif
